`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/05/13 01:13:00
// Design Name: 
// Module Name: ROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ROM(
input wire [6:0]addra,
input wire clka,
output reg [63:0]douta
);

reg [63:0]data[0:127]={
               0,
          456122,
          849611,
         1127499,
         1254653,
         1219187,
         1034284,
          736136,
          378330,
           23545,
         -266158,
         -438949,
         -461259,
         -322989,
          -39087,
          352749,
          797882,
         1233172,
         1596722,
         1837436,
         1922908,
         1844418,
         1618272,
         1283269,
          894694,
          515760,
          207827,
           20909,
          -14067,
          109955,
          375062,
          741142,
         1152081,
         1544437,
         1857255,
         2041483,
         2067568,
         1930020,
         1648268,
         1263660,
          833076,
          420138,
           85383,
         -123094,
         -177060,
          -72507,
          169745,
          507275,
          882633,
         1232235,
         1496210,
         1627669,
         1599968,
         1410850,
         1082801,
          659597,
          199548,
         -233498,
         -580010,
         -793959,
         -849918,
         -746974,
         -508851,
         -180221,
          180221,
          508851,
          746974,
          849918,
          793959,
          580010,
          233498,
         -199548,
         -659597,
        -1082801,
        -1410850,
        -1599968,
        -1627669,
        -1496210,
        -1232235,
         -882633,
         -507275,
         -169745,
           72507,
          177060,
          123094,
          -85383,
         -420138,
         -833076,
        -1263660,
        -1648268,
        -1930020,
        -2067568,
        -2041483,
        -1857255,
        -1544437,
        -1152081,
         -741142,
         -375062,
         -109955,
           14067,
          -20909,
         -207827,
         -515760,
         -894694,
        -1283269,
        -1618272,
        -1844418,
        -1922908,
        -1837436,
        -1596722,
        -1233172,
         -797882,
         -352749,
           39087,
          322989,
          461259,
          438949,
          266158,
          -23545,
         -378330,
         -736136,
        -1034284,
        -1219187,
        -1254653,
        -1127499,
         -849611,
         -456122,
              -0
};

always@(posedge clka)begin
    douta<=data[addra];
end

endmodule
